qweqe:
