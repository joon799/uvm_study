interface counter_if(input logic clk);
    logic rst_n;
    logic en;
    logic [7:0] count;
endinterface

